module not_cell (input wire in,
                output wire out
);
    assign out = ~in;
endmodule